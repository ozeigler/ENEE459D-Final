module testaluregs();
    
endmodule